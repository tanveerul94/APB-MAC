`ifndef OPERAND_WIDTH
  `define OPERAND_WIDTH 8
`endif

`ifndef SLAVE_BASE
	`define	SLAVE_BASE 32'h0000_0000
`endif

interface apb_if(input PCLK);
  bit [31:0] PADDR,PWDATA,PRDATA;
  bit PRESETn,PSELx,PENABLE,PWRITE,PREADY,PSLVERR,BOOTH_READY;
  bit [2*`OPERAND_WIDTH-1:0] BOOTH_OUTPUT;

  modport DRIVER (output PADDR,PWDATA,PRESETn,PSELx,PENABLE,PWRITE,input PCLK,PRDATA,PREADY,PSLVERR,BOOTH_READY);
//  modport MONITOR (input PADDR,PWDATA,PRDATA,PRESETn,PSELx,PENABLE,PWRITE,PREADY,PSLVERR,PCLK);
  modport MONITOR (input PRDATA,PSLVERR,PCLK,BOOTH_OUTPUT);  
    
endinterface 

